`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
// Montek Singh
// 4/12/2017 
//
// PLEASE README!
// ==============
//
// This is a self-checking tester for your full MIPS processor 
// plus memory-mapped IO.
//
// Use this tester carefully!  The names of your top-level input/output
// and internal signals may be different, so modify all of signal names on the
// right-hand-side of the "wire" assigments appearing above the uut
// instantiation.  Observe that the uut itself only has clock and reset inputs
// now, and no debug outputs.  Also, the parameters specifying the names of the
// memory initialization files must match the actual file names.
//
// If you decide not to use some of these internal signals for debugging, you
// may comment the relevant lines out.  Be sure to comment out the
// corresponding "ERROR_*" lines below as well.
//
// Finally, note that in my bitmap memory, each 12-bit color is encoded as
// RRRRGGGGBBBB (i.e., red is most significant).  If you have chosen a different
// order for the red/green/blue color values, you may see ERROR signals for the
// colors light up, but there is no error if you are consistent with your
// RGB ordering.
//
//////////////////////////////////////////////////////////////////////////////////


module project_screentest;

    // Inputs
    logic clk;
    logic reset;

    // Signals inside top-level module uut
    wire [31:0] pc             =uut.pc;                    // PC
    wire [31:0] instr          =uut.instr;                 // instr coming out of instr mem
    wire [31:0] mem_addr       =uut.mem_addr;              // addr sent to data mem
    wire        mem_wr         =uut.mem_wr;                // write enable for data mem
    wire [31:0] mem_readdata   =uut.mem_readdata;          // data read from data mem
    wire [31:0] mem_writedata  =uut.mem_writedata;         // write data for data mem
    
    // Signals inside module uut.mips
    wire        werf           =uut.mips.werf;              // WERF = write enable for register file
    wire  [4:0] alufn          =uut.mips.alufn;             // ALU function
    wire        Z              =uut.mips.Z;                 // Zero flag

    // Signals inside module uut.mips.dp (datapath)
    wire [31:0] ReadData1      =uut.mips.dp.ReadData1;       // Reg[rs]
    wire [31:0] ReadData2      =uut.mips.dp.ReadData2;       // Reg[rt]
    wire [31:0] alu_result     =uut.mips.dp.alu_result;      // ALU's output
    wire [4:0]  reg_writeaddr  =uut.mips.dp.reg_writeaddr;   // destination register
    wire [31:0] reg_writedata  =uut.mips.dp.reg_writedata;   // write data for register file
    wire [31:0] signImm        =uut.mips.dp.signImm;         // sign-/zero-extended immediate
    wire [31:0] aluA           =uut.mips.dp.aluA;            // operand A for ALU
    wire [31:0] aluB           =uut.mips.dp.aluB;            // operand B for ALU

    // Signals inside module uut.mips.c (controller)
    wire [1:0] pcsel           =uut.mips.c.pcsel;
    wire [1:0] wasel           =uut.mips.c.wasel;
    wire sext                  =uut.mips.c.sext;
    wire bsel                  =uut.mips.c.bsel;
    wire [1:0] wdsel           =uut.mips.c.wdsel;
    wire wr                    =uut.mips.c.wr;
    wire [1:0] asel            =uut.mips.c.asel;

    // Signals related to module memIO (memory + memory-mapped IO)
    wire [10:0] smem_addr      =uut.smem_addr;             // address from vgadisplaydriver to access screen mem
    wire [3:0]  charcode       =uut.charcode;              // character code returned by screen mem
    wire dmem_wr               =uut.memIO.dmem_wr;
    wire smem_wr               =uut.memIO.smem_wr;

    // Signals related to module vgadisplaydriver (display driver)
    wire hsync                 =uut.hsync;
    wire vsync                 =uut.vsync;
    wire [3:0] red             =uut.red;
    wire [3:0] green           =uut.green;
    wire [3:0] blue            =uut.blue;
    wire [9:0] x               =uut.display.x;
    wire [9:0] y               =uut.display.y;
    wire [11:0] bmem_addr      =uut.display.bmem_addr;
    wire [11:0] bmem_color     =uut.display.bmem_color;
    

    // Instantiate the Unit Under Test (UUT)
    top uut(
           .clk(clk), 
           .reset(reset)
    );

//
// CHECK ALL VALUES ABOVE THIS LINE
// YOU SHOULD NOT NEED TO MODIFY ANYTHING BELOW
//

    initial begin
        // Initialize Inputs
        clk = 0;
        reset = 0;
   end

   initial begin
      #0.5 clk = 0;
      forever
         #0.5 clk = ~clk;
   end
   
   initial begin
      #200 $finish;
   end
   
   
   
   // SELF-CHECKING CODE
   
   selfcheck_nopause c();

    wire [31:0] c_pc=c.pc;
    wire [31:0] c_instr=c.instr;
    wire [31:0] c_mem_addr=c.mem_addr;
    wire        c_mem_wr=c.mem_wr;
    wire [31:0] c_mem_readdata=c.mem_readdata;
    wire [31:0] c_mem_writedata=c.mem_writedata;
    wire        c_werf=c.werf;
    wire  [4:0] c_alufn=c.alufn;
    wire        c_Z=c.Z;
    wire [31:0] c_ReadData1=c.ReadData1;
    wire [31:0] c_ReadData2=c.ReadData2;
    wire [31:0] c_alu_result=c.alu_result;
    wire [4:0]  c_reg_writeaddr=c.reg_writeaddr;
    wire [31:0] c_reg_writedata=c.reg_writedata;
    wire [31:0] c_signImm=c.signImm;
    wire [31:0] c_aluA=c.aluA;
    wire [31:0] c_aluB=c.aluB;
    wire [1:0]  c_pcsel=c.pcsel;
    wire [1:0]  c_wasel=c.wasel;
    wire        c_sext=c.sext;
    wire        c_bsel=c.bsel;
    wire [1:0]  c_wdsel=c.wdsel;
    wire        c_wr=c.wr;
    wire [1:0]  c_asel=c.asel;
    wire [10:0] c_smem_addr=c.smem_addr;
    wire [3:0]  c_charcode=c.charcode;
    wire        c_dmem_wr=c.dmem_wr;
    wire        c_smem_wr=c.smem_wr;
    wire        c_hsync=c.hsync;
    wire        c_vsync=c.vsync;
    wire [3:0]  c_red=c.red;
    wire [3:0]  c_green=c.green;
    wire [3:0]  c_blue=c.blue;
    wire [9:0]  c_x=c.x;
    wire [9:0]  c_y=c.x;
    wire [11:0] c_bmem_addr=c.bmem_addr;
    wire [11:0] c_bmem_color=c.bmem_color;

  
    function mismatch;  // some trickery needed to match two values with don't cares
        input p, q;      // mismatch in a bit position is ignored if q has an 'x' in that bit
        integer p, q;
        mismatch = (((p ^ q) ^ q) !== q);
    endfunction

    wire ERROR;
    wire ERROR_pc             = mismatch(pc, c.pc) ? 1'bx : 1'b0;
    wire ERROR_instr          = mismatch(instr, c.instr) ? 1'bx : 1'b0;
    wire ERROR_mem_addr       = mismatch(mem_addr, c.mem_addr) ? 1'bx : 1'b0;
    wire ERROR_mem_wr         = mismatch(mem_wr, c.mem_wr) ? 1'bx : 1'b0;
    wire ERROR_mem_readdata   = mismatch(mem_readdata, c.mem_readdata) ? 1'bx : 1'b0;
    wire ERROR_mem_writedata  = c.mem_wr & (mismatch(mem_writedata, c.mem_writedata) ? 1'bx : 1'b0);
    wire ERROR_werf           = mismatch(werf, c.werf) ? 1'bx : 1'b0;
    wire ERROR_alufn          = mismatch(alufn, c.alufn) ? 1'bx : 1'b0;
    wire ERROR_Z              = mismatch(Z, c.Z) ? 1'bx : 1'b0;
    wire ERROR_ReadData1      = mismatch(ReadData1, c.ReadData1) ? 1'bx : 1'b0;
    wire ERROR_ReadData2      = mismatch(ReadData2, c.ReadData2) ? 1'bx : 1'b0;
    wire ERROR_alu_result     = mismatch(alu_result, c.alu_result) ? 1'bx : 1'b0;
    wire ERROR_reg_writeaddr  = c.werf & (mismatch(reg_writeaddr, c.reg_writeaddr) ? 1'bx : 1'b0);
    wire ERROR_reg_writedata  = c.werf & (mismatch(reg_writedata, c.reg_writedata) ? 1'bx : 1'b0);
    wire ERROR_signImm        = mismatch(signImm, c.signImm) ? 1'bx : 1'b0;
    wire ERROR_aluA           = mismatch(aluA, c.aluA) ? 1'bx : 1'b0;
    wire ERROR_aluB           = mismatch(aluB, c.aluB) ? 1'bx : 1'b0;
    wire ERROR_pcsel          = mismatch(pcsel, c.pcsel) ? 1'bx : 1'b0;
    wire ERROR_wasel          = c.werf & (mismatch(wasel, c.wasel) ? 1'bx : 1'b0);
    wire ERROR_sext           = mismatch(sext, c.sext) ? 1'bx : 1'b0;
    wire ERROR_bsel           = mismatch(bsel, c.bsel) ? 1'bx : 1'b0;
    wire ERROR_wdsel          = mismatch(wdsel, c.wdsel) ? 1'bx : 1'b0;
    wire ERROR_wr             = mismatch(wr, c.wr) ? 1'bx : 1'b0;
    wire ERROR_asel           = mismatch(asel, c.asel) ? 1'bx : 1'b0;
    wire ERROR_smem_addr      = mismatch(smem_addr, c.smem_addr) ? 1'bx : 1'b0;
    wire ERROR_charcode       = mismatch(charcode, c.charcode) ? 1'bx : 1'b0;
    wire ERROR_dmem_wr        = mismatch(dmem_wr, c.dmem_wr) ? 1'bx : 1'b0;
    wire ERROR_smem_wr        = mismatch(smem_wr, c.smem_wr) ? 1'bx : 1'b0;
    wire ERROR_hsync          = mismatch(hsync, c.hsync) ? 1'bx : 1'b0;
    wire ERROR_vsync          = mismatch(vsync, c.vsync) ? 1'bx : 1'b0;
    wire ERROR_red            = mismatch(red, c.red) ? 1'bx : 1'b0;
    wire ERROR_green          = mismatch(green, c.green) ? 1'bx : 1'b0;
    wire ERROR_blue           = mismatch(blue, c.blue) ? 1'bx : 1'b0;
    wire ERROR_x              = mismatch(x, c.x) ? 1'bx : 1'b0;
    wire ERROR_y              = mismatch(y, c.y) ? 1'bx : 1'b0;
    wire ERROR_bmem_addr      = mismatch(bmem_addr, c.bmem_addr) ? 1'bx : 1'b0;
    wire ERROR_bmem_color     = mismatch(bmem_color, c.bmem_color) ? 1'bx : 1'b0;

    assign ERROR = ERROR_pc | ERROR_instr | ERROR_mem_addr | ERROR_mem_wr | ERROR_mem_readdata 
              | ERROR_mem_writedata | ERROR_werf | ERROR_alufn | ERROR_Z
              | ERROR_ReadData1 | ERROR_ReadData2 | ERROR_alu_result | ERROR_reg_writeaddr
              | ERROR_reg_writedata | ERROR_signImm | ERROR_aluA | ERROR_aluB
              | ERROR_pcsel | ERROR_wasel | ERROR_sext | ERROR_bsel | ERROR_wdsel | ERROR_wr | ERROR_asel
              | ERROR_smem_addr | ERROR_charcode | ERROR_dmem_wr | ERROR_smem_wr | ERROR_hsync | ERROR_vsync
              | ERROR_red | ERROR_green | ERROR_blue | ERROR_x | ERROR_y | ERROR_bmem_addr | ERROR_bmem_color;


    initial begin
        $monitor("#%02d {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h%h, 32'h%h, 32'h%h, 1'b%b, 32'h%h, 32'h%h, 1'b%b, 5'b%b, 1'b%b, 32'h%h, 32'h%h, 32'h%h, 5'h%h, 32'h%h, 32'h%h, 32'h%h, 32'h%h, 2'b%b, 2'b%b, 1'b%b, 1'b%b, 2'b%b, 1'b%b, 2'b%b};",
                  $time, pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel);
        
        $monitor("#%02d {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h%h, 4'h%h, 1'b%b, 1'b%b, 1'b%b, 1'b%b, 4'h%h, 4'h%h, 4'h%h, 10'h%h, 10'h%h, 12'h%h, 12'h%h};",
                  $time, smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color);
    end
    
endmodule



// CHECKER MODULE

module selfcheck_nopause();
    logic  [31:0] pc;
    logic  [31:0] instr;
    logic  [31:0] mem_addr;
    logic         mem_wr;
    logic  [31:0] mem_readdata;
    logic  [31:0] mem_writedata;
    logic         werf;
    logic   [4:0] alufn;
    logic         Z;
    logic  [31:0] ReadData1;
    logic  [31:0] ReadData2;
    logic  [31:0] alu_result;
    logic  [4:0]  reg_writeaddr;
    logic  [31:0] reg_writedata;
    logic  [31:0] signImm;
    logic  [31:0] aluA;
    logic  [31:0] aluB;
    logic  [1:0] pcsel;
    logic  [1:0] wasel;
    logic        sext;
    logic        bsel;
    logic  [1:0] wdsel;
    logic        wr;
    logic  [1:0] asel;
    logic [10:0] smem_addr;
    logic [3:0]  charcode;
    logic dmem_wr;
    logic smem_wr;
    logic hsync;
    logic vsync;
    logic [3:0] red;
    logic [3:0] green;
    logic [3:0] blue;
    logic [9:0] x;
    logic [9:0] y;
    logic [11:0] bmem_addr;
    logic [11:0] bmem_color;
    
initial begin
fork

#00 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400000, 32'h3c1d1001, 32'h10010000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h10010000, 5'h1d, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#00 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h000, 10'h000, 12'h000, 12'hf00};
#01 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400004, 32'h37bd0100, 32'h10010100, 1'b0, 32'h00000000, 32'h10010000, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'h10010000, 32'h10010100, 5'h1d, 32'h10010100, 32'h00000100, 32'h10010000, 32'h00000100, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#02 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400008, 32'h3c08ffff, 32'hffff0000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'hffff0000, 5'h08, 32'hffff0000, 32'hxxxxffff, 32'h00000010, 32'hxxxxffff, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#03 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040000c, 32'h3508ffff, 32'hffffffff, 1'b0, 32'h00000000, 32'hffff0000, 1'b1, 5'bx0100, 1'b0, 32'hffff0000, 32'hffff0000, 32'hffffffff, 5'h08, 32'hffffffff, 32'h0000ffff, 32'hffff0000, 32'h0000ffff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#04 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400010, 32'h2009ffff, 32'hffffffff, 1'b0, 32'h00000000, 32'hxxxxxxxx, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'hffffffff, 5'h09, 32'hffffffff, 32'hffffffff, 32'h00000000, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#04 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h001, 10'h000, 12'h001, 12'hf00};
#05 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400014, 32'h15090031, 32'h00000000, 1'b0, 32'h00000000, 32'hffffffff, 1'b0, 5'b1xx01, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000031, 32'hffffffff, 32'hffffffff, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#06 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400018, 32'h00084600, 32'hff000000, 1'b0, 32'h00000000, 32'hffffffff, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'hffffffff, 32'hff000000, 5'h08, 32'hff000000, 32'h00004600, 32'h00000018, 32'hffffffff, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#07 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040001c, 32'h3508f000, 32'hff00f000, 1'b0, 32'h00000000, 32'hff000000, 1'b1, 5'bx0100, 1'b0, 32'hff000000, 32'hff000000, 32'hff00f000, 5'h08, 32'hff00f000, 32'h0000f000, 32'hff000000, 32'h0000f000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#08 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400020, 32'h00084203, 32'hffff00f0, 1'b0, 32'h00000000, 32'hff00f000, 1'b1, 5'bx1110, 1'b0, 32'h00000000, 32'hff00f000, 32'hffff00f0, 5'h08, 32'hffff00f0, 32'h00004203, 32'h00000008, 32'hff00f000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#08 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h002, 10'h000, 12'h002, 12'hf00};
#09 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400024, 32'h00084102, 32'h0ffff00f, 1'b0, 32'h00000000, 32'hffff00f0, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'hffff00f0, 32'h0ffff00f, 5'h08, 32'h0ffff00f, 32'h00004102, 32'h00000004, 32'hffff00f0, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#10 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400028, 32'h340a0003, 32'h00000003, 1'b0, 32'h00000000, 32'hxxxxxxxx, 1'b1, 5'bx0100, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000003, 5'h0a, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#11 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040002c, 32'h01495022, 32'h00000004, 1'b0, 32'h00000000, 32'hffffffff, 1'b1, 5'b1xx01, 1'b0, 32'h00000003, 32'hffffffff, 32'h00000004, 5'h0a, 32'h00000004, 32'h00005022, 32'h00000003, 32'hffffffff, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#12 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400030, 32'h01484004, 32'hffff00f0, 1'b0, 32'h00000000, 32'h0ffff00f, 1'b1, 5'bx0010, 1'b0, 32'h00000004, 32'h0ffff00f, 32'hffff00f0, 5'h08, 32'hffff00f0, 32'h00004004, 32'h00000004, 32'h0ffff00f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#12 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h003, 10'h000, 12'h003, 12'hf00};
#13 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400034, 32'h010a582a, 32'h00000001, 1'b0, 32'h00000000, 32'h00000004, 1'b1, 5'b1x011, 1'b0, 32'hffff00f0, 32'h00000004, 32'h00000001, 5'h0b, 32'h00000001, 32'h0000582a, 32'hffff00f0, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#14 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400038, 32'h010a582b, 32'h00000000, 1'b0, 32'h00000000, 32'h00000004, 1'b1, 5'b1x111, 1'b1, 32'hffff00f0, 32'h00000004, 32'h00000000, 5'h0b, 32'h00000000, 32'h0000582b, 32'hffff00f0, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#15 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040003c, 32'h20080005, 32'h00000005, 1'b0, 32'h00000000, 32'hffff00f0, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'hffff00f0, 32'h00000005, 5'h08, 32'h00000005, 32'h00000005, 32'h00000000, 32'h00000005, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#16 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400040, 32'h2d0b000a, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'b1x111, 1'b0, 32'h00000005, 32'h00000000, 32'h00000001, 5'h0b, 32'h00000001, 32'h0000000a, 32'h00000005, 32'h0000000a, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#16 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h004, 10'h000, 12'h004, 12'hf00};
#17 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400044, 32'h2d0b0004, 32'h00000000, 1'b0, 32'h00000000, 32'h00000001, 1'b1, 5'b1x111, 1'b1, 32'h00000005, 32'h00000001, 32'h00000000, 5'h0b, 32'h00000000, 32'h00000004, 32'h00000005, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#18 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400048, 32'h2008fffb, 32'hfffffffb, 1'b0, 32'h00000000, 32'h00000005, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000005, 32'hfffffffb, 5'h08, 32'hfffffffb, 32'hfffffffb, 32'h00000000, 32'hfffffffb, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#19 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040004c, 32'h2d0b0005, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'b1x111, 1'b1, 32'hfffffffb, 32'h00000000, 32'h00000000, 5'h0b, 32'h00000000, 32'h00000005, 32'hfffffffb, 32'h00000005, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#20 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h005, 10'h000, 12'h005, 12'hf00};
#20 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400050, 32'h3c0b1010, 32'h10100000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000000, 32'h10100000, 5'h0b, 32'h10100000, 32'h00001010, 32'h00000010, 32'h00001010, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#21 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400054, 32'h356b1010, 32'h10101010, 1'b0, 32'h00000000, 32'h10100000, 1'b1, 5'bx0100, 1'b0, 32'h10100000, 32'h10100000, 32'h10101010, 5'h0b, 32'h10101010, 32'h00001010, 32'h10100000, 32'h00001010, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#22 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400058, 32'h3c0c0101, 32'h01010000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h01010000, 5'h0c, 32'h01010000, 32'h00000101, 32'h00000010, 32'h00000101, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#23 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040005c, 32'h218c1010, 32'h01011010, 1'b0, 32'hxxxxxxxx, 32'h01010000, 1'b1, 5'b0xx01, 1'b0, 32'h01010000, 32'h01010000, 32'h01011010, 5'h0c, 32'h01011010, 32'h00001010, 32'h01010000, 32'h00001010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#24 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400060, 32'h016c6824, 32'h00001010, 1'b0, 32'h00000000, 32'h01011010, 1'b1, 5'bx0000, 1'b0, 32'h10101010, 32'h01011010, 32'h00001010, 5'h0d, 32'h00001010, 32'h00006824, 32'h10101010, 32'h01011010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#24 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h006, 10'h000, 12'h006, 12'hf00};
#25 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400064, 32'h016c6825, 32'h11111010, 1'b0, 32'hxxxxxxxx, 32'h01011010, 1'b1, 5'bx0100, 1'b0, 32'h10101010, 32'h01011010, 32'h11111010, 5'h0d, 32'h11111010, 32'h00006825, 32'h10101010, 32'h01011010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#26 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400068, 32'h016c6826, 32'h11110000, 1'b0, 32'h00000000, 32'h01011010, 1'b1, 5'bx1000, 1'b0, 32'h10101010, 32'h01011010, 32'h11110000, 5'h0d, 32'h11110000, 32'h00006826, 32'h10101010, 32'h01011010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#27 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040006c, 32'h016c6827, 32'heeeeefef, 1'b0, 32'h00000001, 32'h01011010, 1'b1, 5'bx1100, 1'b0, 32'h10101010, 32'h01011010, 32'heeeeefef, 5'h0d, 32'heeeeefef, 32'h00006827, 32'h10101010, 32'h01011010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#28 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h007, 10'h000, 12'h007, 12'hf00};
#28 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400070, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#29 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400074, 32'h00200821, 32'h10010000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000000, 32'h10010000, 5'h01, 32'h10010000, 32'h00000821, 32'h10010000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#30 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400078, 32'h8c240004, 32'h10010004, 1'b0, 32'h00000003, 32'hxxxxxxxx, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010004, 5'h04, 32'h00000003, 32'h00000004, 32'h10010000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#31 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040007c, 32'h20840002, 32'h00000005, 1'b0, 32'h00000000, 32'h00000003, 1'b1, 5'b0xx01, 1'b0, 32'h00000003, 32'h00000003, 32'h00000005, 5'h04, 32'h00000005, 32'h00000002, 32'h00000003, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#32 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400080, 32'h2484fffe, 32'h00000003, 1'b0, 32'h00000000, 32'h00000005, 1'b1, 5'b0xx01, 1'b0, 32'h00000005, 32'h00000005, 32'h00000003, 5'h04, 32'h00000003, 32'hfffffffe, 32'h00000005, 32'hfffffffe, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#32 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h008, 10'h000, 12'h008, 12'hf00};
#33 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400084, 32'h0c100038, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h00400088, 32'h00000038, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#34 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h23bdfff8, 32'h100100f8, 1'b0, 32'hxxxxxxxx, 32'h10010100, 1'b1, 5'b0xx01, 1'b0, 32'h10010100, 32'h10010100, 32'h100100f8, 5'h1d, 32'h100100f8, 32'hfffffff8, 32'h10010100, 32'hfffffff8, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#35 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'hafbf0004, 32'h100100fc, 1'b1, 32'hxxxxxxxx, 32'h00400088, 1'b0, 5'b0xx01, 1'b0, 32'h100100f8, 32'h00400088, 32'h100100fc, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h100100f8, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#35 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h008, 10'h000, 12'h008, 12'hf00};
#36 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'hafa40000, 32'h100100f8, 1'b1, 32'hxxxxxxxx, 32'h00000003, 1'b0, 5'b0xx01, 1'b0, 32'h100100f8, 32'h00000003, 32'h100100f8, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100100f8, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#36 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h009, 10'h000, 12'h009, 12'hf00};
#37 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h28880002, 32'h00000000, 1'b0, 32'h00000000, 32'hfffffffb, 1'b1, 5'b1x011, 1'b1, 32'h00000003, 32'hfffffffb, 32'h00000000, 5'h08, 32'h00000000, 32'h00000002, 32'h00000003, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#37 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h009, 10'h000, 12'h009, 12'hf00};
#38 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000f0, 32'h11000002, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b0, 5'b1xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#39 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000fc, 32'h2084ffff, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 1'b1, 5'b0xx01, 1'b0, 32'h00000003, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'hffffffff, 32'h00000003, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#40 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400100, 32'h0c100038, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h00400104, 32'h00000038, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#40 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00a, 10'h000, 12'h00a, 12'hf00};
#41 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h23bdfff8, 32'h100100f0, 1'b0, 32'hxxxxxxxx, 32'h100100f8, 1'b1, 5'b0xx01, 1'b0, 32'h100100f8, 32'h100100f8, 32'h100100f0, 5'h1d, 32'h100100f0, 32'hfffffff8, 32'h100100f8, 32'hfffffff8, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#42 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'hafbf0004, 32'h100100f4, 1'b1, 32'hxxxxxxxx, 32'h00400104, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00400104, 32'h100100f4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h100100f0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#42 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00a, 10'h000, 12'h00a, 12'hf00};
#43 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'hafa40000, 32'h100100f0, 1'b1, 32'hxxxxxxxx, 32'h00000002, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000002, 32'h100100f0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100100f0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#44 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h28880002, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'b1x011, 1'b1, 32'h00000002, 32'h00000000, 32'h00000000, 5'h08, 32'h00000000, 32'h00000002, 32'h00000002, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#44 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00b, 10'h000, 12'h00b, 12'hf00};
#45 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000f0, 32'h11000002, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b0, 5'b1xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#46 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000fc, 32'h2084ffff, 32'h00000001, 1'b0, 32'h00000000, 32'h00000002, 1'b1, 5'b0xx01, 1'b0, 32'h00000002, 32'h00000002, 32'h00000001, 5'h04, 32'h00000001, 32'hffffffff, 32'h00000002, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#47 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400100, 32'h0c100038, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h00400104, 32'h00000038, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#48 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h23bdfff8, 32'h100100e8, 1'b0, 32'hxxxxxxxx, 32'h100100f0, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h100100f0, 32'h100100e8, 5'h1d, 32'h100100e8, 32'hfffffff8, 32'h100100f0, 32'hfffffff8, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#48 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00c, 10'h000, 12'h00c, 12'hf00};
#49 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'hafbf0004, 32'h100100ec, 1'b1, 32'hxxxxxxxx, 32'h00400104, 1'b0, 5'b0xx01, 1'b0, 32'h100100e8, 32'h00400104, 32'h100100ec, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h100100e8, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#49 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00c, 10'h000, 12'h00c, 12'hf00};
#50 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'hafa40000, 32'h100100e8, 1'b1, 32'hxxxxxxxx, 32'h00000001, 1'b0, 5'b0xx01, 1'b0, 32'h100100e8, 32'h00000001, 32'h100100e8, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100100e8, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#51 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h28880002, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'b1x011, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'h08, 32'h00000001, 32'h00000002, 32'h00000001, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#51 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00c, 10'h000, 12'h00c, 12'hf00};
#52 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000f0, 32'h11000002, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'h00000002, 32'h00000001, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#52 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00d, 10'h000, 12'h00d, 12'hf00};
#53 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000f4, 32'h00041020, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000001, 32'h00000001, 5'h02, 32'h00000001, 32'h00001020, 32'h00000000, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#54 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000f8, 32'h08100045, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 1'b0, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000045, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#55 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h8fbf0004, 32'h100100ec, 1'b0, 32'h00400104, 32'h00400104, 1'b1, 5'b0xx01, 1'b0, 32'h100100e8, 32'h00400104, 32'h100100ec, 5'h1f, 32'h00400104, 32'h00000004, 32'h100100e8, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#56 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00e, 10'h000, 12'h00e, 12'hf00};
#56 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h23bd0008, 32'h100100f0, 1'b0, 32'h00000002, 32'h100100e8, 1'b1, 5'b0xx01, 1'b0, 32'h100100e8, 32'h100100e8, 32'h100100f0, 5'h1d, 32'h100100f0, 32'h00000008, 32'h100100e8, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#57 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400104, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#58 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'h8fa40000, 32'h100100f0, 1'b0, 32'h00000002, 32'h00000001, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000001, 32'h100100f0, 5'h04, 32'h00000002, 32'h00000000, 32'h100100f0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#59 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'h00441020, 32'h00000003, 1'b0, 32'h00000000, 32'h00000002, 1'b1, 5'b0xx01, 1'b0, 32'h00000001, 32'h00000002, 32'h00000003, 5'h02, 32'h00000003, 32'h00001020, 32'h00000001, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#60 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'h00441020, 32'h00000005, 1'b0, 32'h00000000, 32'h00000002, 1'b1, 5'b0xx01, 1'b0, 32'h00000003, 32'h00000002, 32'h00000005, 5'h02, 32'h00000005, 32'h00001020, 32'h00000003, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#60 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00f, 10'h000, 12'h00f, 12'hf00};
#61 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h2042ffff, 32'h00000004, 1'b0, 32'h00000000, 32'h00000005, 1'b1, 5'b0xx01, 1'b0, 32'h00000005, 32'h00000005, 32'h00000004, 5'h02, 32'h00000004, 32'hffffffff, 32'h00000005, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#62 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h8fbf0004, 32'h100100f4, 1'b0, 32'h00400104, 32'h00400104, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00400104, 32'h100100f4, 5'h1f, 32'h00400104, 32'h00000004, 32'h100100f0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#63 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h23bd0008, 32'h100100f8, 1'b0, 32'h00000003, 32'h100100f0, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h100100f0, 32'h100100f8, 5'h1d, 32'h100100f8, 32'h00000008, 32'h100100f0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#64 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400104, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#64 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h010, 10'h000, 12'h100, 12'h0f0};
#65 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'h8fa40000, 32'h100100f8, 1'b0, 32'h00000003, 32'h00000002, 1'b1, 5'b0xx01, 1'b0, 32'h100100f8, 32'h00000002, 32'h100100f8, 5'h04, 32'h00000003, 32'h00000000, 32'h100100f8, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#66 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'h00441020, 32'h00000007, 1'b0, 32'h00000000, 32'h00000003, 1'b1, 5'b0xx01, 1'b0, 32'h00000004, 32'h00000003, 32'h00000007, 5'h02, 32'h00000007, 32'h00001020, 32'h00000004, 32'h00000003, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#67 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'h00441020, 32'h0000000a, 1'b0, 32'h00000000, 32'h00000003, 1'b1, 5'b0xx01, 1'b0, 32'h00000007, 32'h00000003, 32'h0000000a, 5'h02, 32'h0000000a, 32'h00001020, 32'h00000007, 32'h00000003, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#68 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h2042ffff, 32'h00000009, 1'b0, 32'h00000000, 32'h0000000a, 1'b1, 5'b0xx01, 1'b0, 32'h0000000a, 32'h0000000a, 32'h00000009, 5'h02, 32'h00000009, 32'hffffffff, 32'h0000000a, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#68 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h011, 10'h000, 12'h101, 12'h0f0};
#69 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h8fbf0004, 32'h100100fc, 1'b0, 32'h00400088, 32'h00400104, 1'b1, 5'b0xx01, 1'b0, 32'h100100f8, 32'h00400104, 32'h100100fc, 5'h1f, 32'h00400088, 32'h00000004, 32'h100100f8, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#70 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h23bd0008, 32'h10010100, 1'b0, 32'h00000000, 32'h100100f8, 1'b1, 5'b0xx01, 1'b0, 32'h100100f8, 32'h100100f8, 32'h10010100, 5'h1d, 32'h10010100, 32'h00000008, 32'h100100f8, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#71 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400088, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#72 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h012, 10'h000, 12'h102, 12'h0f0};
#72 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400088, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#73 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040008c, 32'h00200821, 32'h10010000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000000, 32'h10010000, 5'h01, 32'h10010000, 32'h00000821, 32'h10010000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#74 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400090, 32'hac220000, 32'h10010000, 1'b1, 32'h00000000, 32'h00000009, 1'b0, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000009, 32'h10010000, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010000, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#74 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h012, 10'h000, 12'h102, 12'h0f0};
#75 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400094, 32'h200403e8, 32'h000003e8, 1'b0, 32'h00000000, 32'h00000003, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h000003e8, 5'h04, 32'h000003e8, 32'h000003e8, 32'h00000000, 32'h000003e8, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#75 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h012, 10'h000, 12'h102, 12'h0f0};
#76 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400098, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#76 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h013, 10'h000, 12'h103, 12'h0f0};
#77 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040009c, 32'h24050000, 32'h00000000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 5'h05, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#78 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000a0, 32'h24060000, 32'h00000000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 5'h06, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#79 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000a4, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h000003e8, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h000003e8, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#80 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000a8, 32'h0c100053, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h004000ac, 32'h00000053, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#80 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h014, 10'h000, 12'h104, 12'h0f0};
#81 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040014c, 32'h23bdfff0, 32'h100100f0, 1'b0, 32'h00000002, 32'h10010100, 1'b1, 5'b0xx01, 1'b0, 32'h10010100, 32'h10010100, 32'h100100f0, 5'h1d, 32'h100100f0, 32'hfffffff0, 32'h10010100, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#82 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400150, 32'hafbf000c, 32'h100100fc, 1'b1, 32'h00400088, 32'h004000ac, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h004000ac, 32'h100100fc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h100100f0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#82 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h014, 10'h000, 12'h104, 12'h0f0};
#83 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400154, 32'hafa80008, 32'h100100f8, 1'b1, 32'h00000003, 32'h00000001, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000001, 32'h100100f8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h100100f0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#84 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400158, 32'hafa90004, 32'h100100f4, 1'b1, 32'h00400104, 32'hffffffff, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'hffffffff, 32'h100100f4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h100100f0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#84 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h015, 10'h000, 12'h105, 12'h0f0};
#85 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040015c, 32'hafaa0000, 32'h100100f0, 1'b1, 32'h00000002, 32'h00000004, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000004, 32'h100100f0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100100f0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#86 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400160, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000000, 32'h10010000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#86 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h015, 10'h000, 12'h105, 12'h0f0};
#87 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400164, 32'h34280000, 32'h10020000, 1'b0, 32'h00000000, 32'h00000001, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#88 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400168, 32'h00064940, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004940, 32'h00000005, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#88 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h016, 10'h000, 12'h106, 12'h0f0};
#89 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040016c, 32'h000650c0, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h0a, 32'h00000000, 32'h000050c0, 32'h00000003, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#90 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h012a4820, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004820, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#91 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'h01254820, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004820, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#92 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h017, 10'h000, 12'h107, 12'h0f0};
#92 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'h00094880, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004880, 32'h00000002, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#93 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'h01094020, 32'h10020000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000000, 32'h10020000, 5'h08, 32'h10020000, 32'h00004020, 32'h10020000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#94 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'had040000, 32'h10020000, 1'b1, 32'h00000000, 32'h00000002, 1'b0, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000002, 32'h10020000, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#94 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h017, 10'h000, 12'h107, 12'h0f0};
#95 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h8fbf000c, 32'h100100fc, 1'b0, 32'h004000ac, 32'h004000ac, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h004000ac, 32'h100100fc, 5'h1f, 32'h004000ac, 32'h0000000c, 32'h100100f0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#95 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h017, 10'h000, 12'h107, 12'h0f0};
#96 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h018, 10'h000, 12'h108, 12'h0f0};
#96 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h8fa80008, 32'h100100f8, 1'b0, 32'h00000001, 32'h10020000, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h10020000, 32'h100100f8, 5'h08, 32'h00000001, 32'h00000008, 32'h100100f0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#97 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h8fa90004, 32'h100100f4, 1'b0, 32'hffffffff, 32'h00000000, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000000, 32'h100100f4, 5'h09, 32'hffffffff, 32'h00000004, 32'h100100f0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#98 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h8faa0000, 32'h100100f0, 1'b0, 32'h00000004, 32'h00000000, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000000, 32'h100100f0, 5'h0a, 32'h00000004, 32'h00000000, 32'h100100f0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#99 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h23bd0010, 32'h10010100, 1'b0, 32'h00000009, 32'h100100f0, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h100100f0, 32'h10010100, 5'h1d, 32'h10010100, 32'h00000010, 32'h100100f0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#100 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000ac, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#100 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h019, 10'h000, 12'h109, 12'h0f0};
#101 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000ac, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#102 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000b0, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#103 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000b4, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#104 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000b8, 32'h0c100053, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h004000bc, 32'h00000053, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#104 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01a, 10'h000, 12'h10a, 12'h0f0};
#105 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040014c, 32'h23bdfff0, 32'h100100f0, 1'b0, 32'h00000004, 32'h10010100, 1'b1, 5'b0xx01, 1'b0, 32'h10010100, 32'h10010100, 32'h100100f0, 5'h1d, 32'h100100f0, 32'hfffffff0, 32'h10010100, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#106 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400150, 32'hafbf000c, 32'h100100fc, 1'b1, 32'h004000ac, 32'h004000bc, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h004000bc, 32'h100100fc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h100100f0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#106 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01a, 10'h000, 12'h10a, 12'h0f0};
#107 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400154, 32'hafa80008, 32'h100100f8, 1'b1, 32'h00000001, 32'h00000001, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000001, 32'h100100f8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h100100f0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#108 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01b, 10'h000, 12'h10b, 12'h0f0};
#108 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400158, 32'hafa90004, 32'h100100f4, 1'b1, 32'hffffffff, 32'hffffffff, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'hffffffff, 32'h100100f4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h100100f0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#109 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040015c, 32'hafaa0000, 32'h100100f0, 1'b1, 32'h00000004, 32'h00000004, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000004, 32'h100100f0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100100f0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#110 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400160, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000002, 32'h10020000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#110 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01b, 10'h000, 12'h10b, 12'h0f0};
#111 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400164, 32'h34280000, 32'h10020000, 1'b0, 32'h00000002, 32'h00000001, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#112 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400168, 32'h00064940, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004940, 32'h00000005, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#112 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01c, 10'h000, 12'h10c, 12'h0f0};
#113 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040016c, 32'h000650c0, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h0a, 32'h00000000, 32'h000050c0, 32'h00000003, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#114 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h012a4820, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004820, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#115 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'h01254820, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004820, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#116 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01d, 10'h000, 12'h10d, 12'h0f0};
#116 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'h00094880, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004880, 32'h00000002, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#117 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'h01094020, 32'h10020000, 1'b0, 32'h00000002, 32'h00000000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000000, 32'h10020000, 5'h08, 32'h10020000, 32'h00004020, 32'h10020000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#118 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'had040000, 32'h10020000, 1'b1, 32'h00000002, 32'h00000003, 1'b0, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000003, 32'h10020000, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#118 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01d, 10'h000, 12'h10d, 12'h0f0};
#119 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h8fbf000c, 32'h100100fc, 1'b0, 32'h004000bc, 32'h004000bc, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h004000bc, 32'h100100fc, 5'h1f, 32'h004000bc, 32'h0000000c, 32'h100100f0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#119 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01d, 10'h000, 12'h10d, 12'h0f0};
#120 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01e, 10'h000, 12'h10e, 12'h0f0};
#120 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h8fa80008, 32'h100100f8, 1'b0, 32'h00000001, 32'h10020000, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h10020000, 32'h100100f8, 5'h08, 32'h00000001, 32'h00000008, 32'h100100f0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#121 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h8fa90004, 32'h100100f4, 1'b0, 32'hffffffff, 32'h00000000, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000000, 32'h100100f4, 5'h09, 32'hffffffff, 32'h00000004, 32'h100100f0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#122 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h8faa0000, 32'h100100f0, 1'b0, 32'h00000004, 32'h00000000, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000000, 32'h100100f0, 5'h0a, 32'h00000004, 32'h00000000, 32'h100100f0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#123 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h23bd0010, 32'h10010100, 1'b0, 32'h00000009, 32'h100100f0, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h100100f0, 32'h10010100, 5'h1d, 32'h10010100, 32'h00000010, 32'h100100f0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#124 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000bc, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#124 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01f, 10'h000, 12'h10f, 12'h0f0};
#125 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000bc, 32'h20a50001, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000000, 32'h00000001, 5'h05, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#126 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000c0, 32'h20c60001, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000000, 32'h00000001, 5'h06, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#127 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000c4, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 1'b1, 5'b1x011, 1'b0, 32'h00000001, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000001, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#128 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h020, 10'h000, 12'h000, 12'hf00};
#128 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#129 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000a4, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#130 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000a8, 32'h0c100053, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h004000ac, 32'h00000053, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#131 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040014c, 32'h23bdfff0, 32'h100100f0, 1'b0, 32'h00000004, 32'h10010100, 1'b1, 5'b0xx01, 1'b0, 32'h10010100, 32'h10010100, 32'h100100f0, 5'h1d, 32'h100100f0, 32'hfffffff0, 32'h10010100, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#132 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400150, 32'hafbf000c, 32'h100100fc, 1'b1, 32'h004000bc, 32'h004000ac, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h004000ac, 32'h100100fc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h100100f0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#132 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h021, 10'h000, 12'h001, 12'hf00};
#133 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400154, 32'hafa80008, 32'h100100f8, 1'b1, 32'h00000001, 32'h00000001, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000001, 32'h100100f8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h100100f0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#134 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400158, 32'hafa90004, 32'h100100f4, 1'b1, 32'hffffffff, 32'hffffffff, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'hffffffff, 32'h100100f4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h100100f0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#135 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040015c, 32'hafaa0000, 32'h100100f0, 1'b1, 32'h00000004, 32'h00000004, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000004, 32'h100100f0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100100f0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#136 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h022, 10'h000, 12'h002, 12'hf00};
#136 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400160, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#137 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400164, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#138 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400168, 32'h00064940, 32'h00000020, 1'b0, 32'h00000000, 32'h00000001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h00000020, 5'h09, 32'h00000020, 32'h00004940, 32'h00000005, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#139 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040016c, 32'h000650c0, 32'h00000008, 1'b0, 32'h00000000, 32'h00000001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h00000008, 5'h0a, 32'h00000008, 32'h000050c0, 32'h00000003, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#140 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h023, 10'h000, 12'h003, 12'hf00};
#140 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h012a4820, 32'h00000028, 1'b0, 32'h00000000, 32'h00000008, 1'b1, 5'b0xx01, 1'b0, 32'h00000020, 32'h00000008, 32'h00000028, 5'h09, 32'h00000028, 32'h00004820, 32'h00000020, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#141 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'h01254820, 32'h00000029, 1'b0, 32'h00000000, 32'h00000001, 1'b1, 5'b0xx01, 1'b0, 32'h00000028, 32'h00000001, 32'h00000029, 5'h09, 32'h00000029, 32'h00004820, 32'h00000028, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#142 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'h00094880, 32'h000000a4, 1'b0, 32'h00000000, 32'h00000029, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000029, 32'h000000a4, 5'h09, 32'h000000a4, 32'h00004880, 32'h00000002, 32'h00000029, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#143 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'h01094020, 32'h100200a4, 1'b0, 32'h00000001, 32'h000000a4, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000000a4, 32'h100200a4, 5'h08, 32'h100200a4, 32'h00004020, 32'h10020000, 32'h000000a4, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#144 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'had040000, 32'h100200a4, 1'b1, 32'h00000001, 32'h00000002, 1'b0, 5'b0xx01, 1'b0, 32'h100200a4, 32'h00000002, 32'h100200a4, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100200a4, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#144 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h024, 10'h000, 12'h004, 12'hf00};
#145 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h8fbf000c, 32'h100100fc, 1'b0, 32'h004000ac, 32'h004000ac, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h004000ac, 32'h100100fc, 5'h1f, 32'h004000ac, 32'h0000000c, 32'h100100f0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#145 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h024, 10'h000, 12'h004, 12'hf00};
#146 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h8fa80008, 32'h100100f8, 1'b0, 32'h00000001, 32'h100200a4, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h100200a4, 32'h100100f8, 5'h08, 32'h00000001, 32'h00000008, 32'h100100f0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#147 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h8fa90004, 32'h100100f4, 1'b0, 32'hffffffff, 32'h000000a4, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h000000a4, 32'h100100f4, 5'h09, 32'hffffffff, 32'h00000004, 32'h100100f0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#148 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h8faa0000, 32'h100100f0, 1'b0, 32'h00000004, 32'h00000008, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000008, 32'h100100f0, 5'h0a, 32'h00000004, 32'h00000000, 32'h100100f0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#148 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h025, 10'h000, 12'h005, 12'hf00};
#149 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h23bd0010, 32'h10010100, 1'b0, 32'h00000009, 32'h100100f0, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h100100f0, 32'h10010100, 5'h1d, 32'h10010100, 32'h00000010, 32'h100100f0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#150 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000ac, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#151 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000ac, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#152 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000b0, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#152 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h026, 10'h000, 12'h006, 12'hf00};
#153 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000b4, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#154 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000b8, 32'h0c100053, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h004000bc, 32'h00000053, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#155 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040014c, 32'h23bdfff0, 32'h100100f0, 1'b0, 32'h00000004, 32'h10010100, 1'b1, 5'b0xx01, 1'b0, 32'h10010100, 32'h10010100, 32'h100100f0, 5'h1d, 32'h100100f0, 32'hfffffff0, 32'h10010100, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#156 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400150, 32'hafbf000c, 32'h100100fc, 1'b1, 32'h004000ac, 32'h004000bc, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h004000bc, 32'h100100fc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h100100f0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#156 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h027, 10'h000, 12'h007, 12'hf00};
#157 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400154, 32'hafa80008, 32'h100100f8, 1'b1, 32'h00000001, 32'h00000001, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000001, 32'h100100f8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h100100f0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#158 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400158, 32'hafa90004, 32'h100100f4, 1'b1, 32'hffffffff, 32'hffffffff, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'hffffffff, 32'h100100f4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h100100f0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#159 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040015c, 32'hafaa0000, 32'h100100f0, 1'b1, 32'h00000004, 32'h00000004, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000004, 32'h100100f0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100100f0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#160 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h028, 10'h000, 12'h008, 12'hf00};
#160 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400160, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#161 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400164, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#162 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400168, 32'h00064940, 32'h00000020, 1'b0, 32'h00000000, 32'h00000001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h00000020, 5'h09, 32'h00000020, 32'h00004940, 32'h00000005, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#163 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040016c, 32'h000650c0, 32'h00000008, 1'b0, 32'h00000000, 32'h00000001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h00000008, 5'h0a, 32'h00000008, 32'h000050c0, 32'h00000003, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#164 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h029, 10'h000, 12'h009, 12'hf00};
#164 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h012a4820, 32'h00000028, 1'b0, 32'h00000000, 32'h00000008, 1'b1, 5'b0xx01, 1'b0, 32'h00000020, 32'h00000008, 32'h00000028, 5'h09, 32'h00000028, 32'h00004820, 32'h00000020, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#165 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'h01254820, 32'h00000029, 1'b0, 32'h00000000, 32'h00000001, 1'b1, 5'b0xx01, 1'b0, 32'h00000028, 32'h00000001, 32'h00000029, 5'h09, 32'h00000029, 32'h00004820, 32'h00000028, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#166 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'h00094880, 32'h000000a4, 1'b0, 32'h00000000, 32'h00000029, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000029, 32'h000000a4, 5'h09, 32'h000000a4, 32'h00004880, 32'h00000002, 32'h00000029, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#167 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'h01094020, 32'h100200a4, 1'b0, 32'h00000002, 32'h000000a4, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000000a4, 32'h100200a4, 5'h08, 32'h100200a4, 32'h00004020, 32'h10020000, 32'h000000a4, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#168 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'had040000, 32'h100200a4, 1'b1, 32'h00000002, 32'h00000003, 1'b0, 5'b0xx01, 1'b0, 32'h100200a4, 32'h00000003, 32'h100200a4, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100200a4, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#168 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02a, 10'h000, 12'h00a, 12'hf00};
#169 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h8fbf000c, 32'h100100fc, 1'b0, 32'h004000bc, 32'h004000bc, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h004000bc, 32'h100100fc, 5'h1f, 32'h004000bc, 32'h0000000c, 32'h100100f0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#169 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02a, 10'h000, 12'h00a, 12'hf00};
#170 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h8fa80008, 32'h100100f8, 1'b0, 32'h00000001, 32'h100200a4, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h100200a4, 32'h100100f8, 5'h08, 32'h00000001, 32'h00000008, 32'h100100f0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#171 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h8fa90004, 32'h100100f4, 1'b0, 32'hffffffff, 32'h000000a4, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h000000a4, 32'h100100f4, 5'h09, 32'hffffffff, 32'h00000004, 32'h100100f0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#172 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h8faa0000, 32'h100100f0, 1'b0, 32'h00000004, 32'h00000008, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000008, 32'h100100f0, 5'h0a, 32'h00000004, 32'h00000000, 32'h100100f0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#172 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02b, 10'h000, 12'h00b, 12'hf00};
#173 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h23bd0010, 32'h10010100, 1'b0, 32'h00000009, 32'h100100f0, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h100100f0, 32'h10010100, 5'h1d, 32'h10010100, 32'h00000010, 32'h100100f0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#174 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000bc, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#175 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000bc, 32'h20a50001, 32'h00000002, 1'b0, 32'h00000000, 32'h00000001, 1'b1, 5'b0xx01, 1'b0, 32'h00000001, 32'h00000001, 32'h00000002, 5'h05, 32'h00000002, 32'h00000001, 32'h00000001, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#176 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000c0, 32'h20c60001, 32'h00000002, 1'b0, 32'h00000000, 32'h00000001, 1'b1, 5'b0xx01, 1'b0, 32'h00000001, 32'h00000001, 32'h00000002, 5'h06, 32'h00000002, 32'h00000001, 32'h00000001, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#176 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02c, 10'h000, 12'h00c, 12'hf00};
#177 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000c4, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 1'b1, 5'b1x011, 1'b0, 32'h00000002, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000002, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#178 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#179 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000a4, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#180 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h004000a8, 32'h0c100053, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h004000ac, 32'h00000053, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#180 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02d, 10'h000, 12'h00d, 12'hf00};
#181 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040014c, 32'h23bdfff0, 32'h100100f0, 1'b0, 32'h00000004, 32'h10010100, 1'b1, 5'b0xx01, 1'b0, 32'h10010100, 32'h10010100, 32'h100100f0, 5'h1d, 32'h100100f0, 32'hfffffff0, 32'h10010100, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#182 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400150, 32'hafbf000c, 32'h100100fc, 1'b1, 32'h004000bc, 32'h004000ac, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h004000ac, 32'h100100fc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h100100f0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#182 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02d, 10'h000, 12'h00d, 12'hf00};
#183 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400154, 32'hafa80008, 32'h100100f8, 1'b1, 32'h00000001, 32'h00000001, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000001, 32'h100100f8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h100100f0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#184 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02e, 10'h000, 12'h00e, 12'hf00};
#184 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400158, 32'hafa90004, 32'h100100f4, 1'b1, 32'hffffffff, 32'hffffffff, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'hffffffff, 32'h100100f4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h100100f0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#185 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040015c, 32'hafaa0000, 32'h100100f0, 1'b1, 32'h00000004, 32'h00000004, 1'b0, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000004, 32'h100100f0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100100f0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#186 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400160, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#186 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02e, 10'h000, 12'h00e, 12'hf00};
#187 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400164, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#188 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400168, 32'h00064940, 32'h00000040, 1'b0, 32'h00000000, 32'h00000002, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000002, 32'h00000040, 5'h09, 32'h00000040, 32'h00004940, 32'h00000005, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#188 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02f, 10'h000, 12'h00f, 12'hf00};
#189 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040016c, 32'h000650c0, 32'h00000010, 1'b0, 32'h00000000, 32'h00000002, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000002, 32'h00000010, 5'h0a, 32'h00000010, 32'h000050c0, 32'h00000003, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#190 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h012a4820, 32'h00000050, 1'b0, 32'h00000000, 32'h00000010, 1'b1, 5'b0xx01, 1'b0, 32'h00000040, 32'h00000010, 32'h00000050, 5'h09, 32'h00000050, 32'h00004820, 32'h00000040, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#191 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'h01254820, 32'h00000052, 1'b0, 32'h00000000, 32'h00000002, 1'b1, 5'b0xx01, 1'b0, 32'h00000050, 32'h00000002, 32'h00000052, 5'h09, 32'h00000052, 32'h00004820, 32'h00000050, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#192 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'h00094880, 32'h00000148, 1'b0, 32'h00000000, 32'h00000052, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000052, 32'h00000148, 5'h09, 32'h00000148, 32'h00004880, 32'h00000002, 32'h00000052, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#192 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h030, 10'h000, 12'h100, 12'h0f0};
#193 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'h01094020, 32'h10020148, 1'b0, 32'h00000000, 32'h00000148, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000148, 32'h10020148, 5'h08, 32'h10020148, 32'h00004020, 32'h10020000, 32'h00000148, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#194 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'had040000, 32'h10020148, 1'b1, 32'h00000000, 32'h00000002, 1'b0, 5'b0xx01, 1'b0, 32'h10020148, 32'h00000002, 32'h10020148, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020148, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#194 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h030, 10'h000, 12'h100, 12'h0f0};
#195 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h8fbf000c, 32'h100100fc, 1'b0, 32'h004000ac, 32'h004000ac, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h004000ac, 32'h100100fc, 5'h1f, 32'h004000ac, 32'h0000000c, 32'h100100f0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#195 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h030, 10'h000, 12'h100, 12'h0f0};
#196 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h031, 10'h000, 12'h101, 12'h0f0};
#196 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h8fa80008, 32'h100100f8, 1'b0, 32'h00000001, 32'h10020148, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h10020148, 32'h100100f8, 5'h08, 32'h00000001, 32'h00000008, 32'h100100f0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#197 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h8fa90004, 32'h100100f4, 1'b0, 32'hffffffff, 32'h00000148, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000148, 32'h100100f4, 5'h09, 32'hffffffff, 32'h00000004, 32'h100100f0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#198 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h8faa0000, 32'h100100f0, 1'b0, 32'h00000004, 32'h00000010, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h00000010, 32'h100100f0, 5'h0a, 32'h00000004, 32'h00000000, 32'h100100f0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#199 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h23bd0010, 32'h10010100, 1'b0, 32'h00000009, 32'h100100f0, 1'b1, 5'b0xx01, 1'b0, 32'h100100f0, 32'h100100f0, 32'h10010100, 5'h1d, 32'h10010100, 32'h00000010, 32'h100100f0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};

join
end

endmodule
